module Digital_Equalizer(
	clk,
	clk_for_fir,
	rst_n,
	fir_ready,
	in,
	//tap_f0,tap_f1,tap_f2,tap_f3,tap_f4,tap_f5,tap_f6,tap_f7,
	gain,
	out,
	);
		
	input clk;
	input clk_for_fir;
	input rst_n;
	input fir_ready;
	input signed [15:0] in;
	//input signed [79:0] tap_f0,tap_f1,tap_f2,tap_f3,tap_f4,tap_f5,tap_f6,tap_f7;
	input signed [39:0] gain;
	output signed [15:0] out;
	
	wire signed [239:0] tap_f1,tap_f2,tap_f3,tap_f4,tap_f5,tap_f6,tap_f7,tap_f8;
	
	wire signed [31:0] fir_out1,fir_out2,fir_out3,fir_out4,fir_out5,fir_out6,fir_out7,fir_out8;
	wire signed [20:0] gain_out1,gain_out2,gain_out3,gain_out4,gain_out5,gain_out6,gain_out7,gain_out8;
		
	assign	tap_f1=240'b000000010101001100000010000101100000010000111000000001110100111100001010101111110000110111011010000100000000001000010000110010000001000000000101000011011101111100001010110001010000011101010101000001000011110100000010000110000000000101010011;
	assign	tap_f2=240'b111111111110111011111111111011011111111111101000111111111110110111111111111111100000000000010100000000000010100000000000001100000000000000101000000000000001010011111111111111101111111111101101111111111110100011111111111011001111111111101110;
	assign	tap_f3=240'b111111110110010111111111010011101111111100011001111111110011100111111111110101000000000010111010000000011000010100000001110101100000000110000110000000001011101011111111110101001111111100111000111111110001011111111111010011011111111101100101;
	assign	tap_f4=240'b111111101111001111111110010110011111110100110110111111001110001011111110011110010000000111000100000001010001111100000110100010010000010100100000000000011100010111111110011110001111110011011111111111010011001111111110010101111111111011110011;
	assign	tap_f5=240'b000000001010101000000000000001001111110110010000111110011000101111111000101010111111111100001100000010010101001000001110011010010000100101010100111111110000101111111000101001111111100110000110111111011000110100000000000001000000000010101010;
	assign	tap_f6=240'b111111110100011100000000010101000000010000010100000000110001110011110101100011001111000010001110000001101110001000011000011100010000011011100011111100001000100011110101100001100000001100011111000001000001100100000000010101011111111101000111;
	assign	tap_f7=240'b000000001010010011111111011001111111111111010101111110111001000100010000110100001111010000001100111001111110010100101111101001011110011111100001111101000000100000010000110110011111101110001101111111111101010011111111011001100000000010100100;
	assign	tap_f8=240'b000000000000000000000000000101111111111101010010000000100110100111111010001111100000101001001000111100011010011100010000000000101111000110100111000010100100100011111010001111100000001001101001111111110101001000000000000101110000000000000000;


	fir_v2 F1 (clk_for_fir,rst_n,fir_ready,in,tap_f1,fir_out1);
	fir_v2 F2 (clk_for_fir,rst_n,fir_ready,in,tap_f2,fir_out2);
	fir_v2 F3 (clk_for_fir,rst_n,fir_ready,in,tap_f3,fir_out3);
	fir_v2 F4 (clk_for_fir,rst_n,fir_ready,in,tap_f4,fir_out4);
	fir_v2 F5 (clk_for_fir,rst_n,fir_ready,in,tap_f5,fir_out5);
	fir_v2 F6 (clk_for_fir,rst_n,fir_ready,in,tap_f6,fir_out6);
	fir_v2 F7 (clk_for_fir,rst_n,fir_ready,in,tap_f7,fir_out7);
	fir_v2 F8 (clk_for_fir,rst_n,fir_ready,in,tap_f8,fir_out8);
	
	slider_gain G1 (clk,rst_n,fir_out1[31:16],gain[4:0],gain_out1);
	slider_gain G2 (clk,rst_n,fir_out2[31:16],gain[9:5],gain_out2);
	slider_gain G3 (clk,rst_n,fir_out3[31:16],gain[14:10],gain_out3);
	slider_gain G4 (clk,rst_n,fir_out4[31:16],gain[19:15],gain_out4);
	slider_gain G5 (clk,rst_n,fir_out5[31:16],gain[24:20],gain_out5);
	slider_gain G6 (clk,rst_n,fir_out6[31:16],gain[29:25],gain_out6);
	slider_gain G7 (clk,rst_n,fir_out7[31:16],gain[34:30],gain_out7);
	slider_gain G8 (clk,rst_n,fir_out8[31:16],gain[39:35],gain_out8);
	
	add_data A (clk,rst_n,{gain_out1,gain_out2,gain_out3,gain_out4,gain_out5,gain_out6,gain_out7,gain_out8},out);
	

endmodule
	